library verilog;
use verilog.vl_types.all;
entity Decoder_5_to_32_vlg_vec_tst is
end Decoder_5_to_32_vlg_vec_tst;
