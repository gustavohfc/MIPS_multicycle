library verilog;
use verilog.vl_types.all;
entity Coprocessador_Arithmetic_Unit_vlg_vec_tst is
end Coprocessador_Arithmetic_Unit_vlg_vec_tst;
