library verilog;
use verilog.vl_types.all;
entity Shift_right_arithmetic_vlg_vec_tst is
end Shift_right_arithmetic_vlg_vec_tst;
