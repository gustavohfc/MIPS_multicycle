library verilog;
use verilog.vl_types.all;
entity Controle_ALU_vlg_vec_tst is
end Controle_ALU_vlg_vec_tst;
