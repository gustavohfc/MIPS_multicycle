library verilog;
use verilog.vl_types.all;
entity Extensao_de_sinal_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end Extensao_de_sinal_vlg_check_tst;
