library verilog;
use verilog.vl_types.all;
entity Instruction_register_vlg_vec_tst is
end Instruction_register_vlg_vec_tst;
