library verilog;
use verilog.vl_types.all;
entity Extensao_de_sinal_vlg_vec_tst is
end Extensao_de_sinal_vlg_vec_tst;
