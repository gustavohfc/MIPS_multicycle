library verilog;
use verilog.vl_types.all;
entity lpm_constant0 is
    port(
        result          : out    vl_logic_vector(4 downto 0)
    );
end lpm_constant0;
