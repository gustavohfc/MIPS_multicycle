library verilog;
use verilog.vl_types.all;
entity Decoder_5_to_32_vlg_check_tst is
    port(
        out_0           : in     vl_logic;
        out_1           : in     vl_logic;
        out_2           : in     vl_logic;
        out_3           : in     vl_logic;
        out_4           : in     vl_logic;
        out_5           : in     vl_logic;
        out_6           : in     vl_logic;
        out_7           : in     vl_logic;
        out_8           : in     vl_logic;
        out_9           : in     vl_logic;
        out_10          : in     vl_logic;
        out_11          : in     vl_logic;
        out_12          : in     vl_logic;
        out_13          : in     vl_logic;
        out_14          : in     vl_logic;
        out_15          : in     vl_logic;
        out_16          : in     vl_logic;
        out_17          : in     vl_logic;
        out_18          : in     vl_logic;
        out_19          : in     vl_logic;
        out_20          : in     vl_logic;
        out_21          : in     vl_logic;
        out_22          : in     vl_logic;
        out_23          : in     vl_logic;
        out_24          : in     vl_logic;
        out_25          : in     vl_logic;
        out_26          : in     vl_logic;
        out_27          : in     vl_logic;
        out_28          : in     vl_logic;
        out_29          : in     vl_logic;
        out_30          : in     vl_logic;
        out_31          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Decoder_5_to_32_vlg_check_tst;
