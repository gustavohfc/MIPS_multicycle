library verilog;
use verilog.vl_types.all;
entity Coprocessador_vlg_vec_tst is
end Coprocessador_vlg_vec_tst;
