library verilog;
use verilog.vl_types.all;
entity word_register_vlg_vec_tst is
end word_register_vlg_vec_tst;
