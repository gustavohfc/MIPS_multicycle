library verilog;
use verilog.vl_types.all;
entity Decoder_5_to_32 is
    port(
        out_0           : out    vl_logic;
        RegNumber       : in     vl_logic_vector(4 downto 0);
        out_1           : out    vl_logic;
        out_2           : out    vl_logic;
        out_3           : out    vl_logic;
        out_4           : out    vl_logic;
        out_5           : out    vl_logic;
        out_6           : out    vl_logic;
        out_7           : out    vl_logic;
        out_8           : out    vl_logic;
        out_9           : out    vl_logic;
        out_10          : out    vl_logic;
        out_11          : out    vl_logic;
        out_12          : out    vl_logic;
        out_13          : out    vl_logic;
        out_14          : out    vl_logic;
        out_15          : out    vl_logic;
        out_16          : out    vl_logic;
        out_17          : out    vl_logic;
        out_18          : out    vl_logic;
        out_19          : out    vl_logic;
        out_20          : out    vl_logic;
        out_21          : out    vl_logic;
        out_22          : out    vl_logic;
        out_23          : out    vl_logic;
        out_24          : out    vl_logic;
        out_25          : out    vl_logic;
        out_26          : out    vl_logic;
        out_27          : out    vl_logic;
        out_28          : out    vl_logic;
        out_29          : out    vl_logic;
        out_30          : out    vl_logic;
        out_31          : out    vl_logic
    );
end Decoder_5_to_32;
