library verilog;
use verilog.vl_types.all;
entity lpm_constant1 is
    port(
        result          : out    vl_logic_vector(31 downto 0)
    );
end lpm_constant1;
