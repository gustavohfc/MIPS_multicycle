library verilog;
use verilog.vl_types.all;
entity lpm_constant2_lpm_constant_c19 is
    port(
        result          : out    vl_logic_vector(31 downto 0)
    );
end lpm_constant2_lpm_constant_c19;
