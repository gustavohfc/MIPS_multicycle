library verilog;
use verilog.vl_types.all;
entity Banco_de_registradores_vlg_vec_tst is
end Banco_de_registradores_vlg_vec_tst;
