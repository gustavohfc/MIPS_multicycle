library verilog;
use verilog.vl_types.all;
entity RAM is
    port(
        address         : in     vl_logic_vector(13 downto 0);
        data            : in     vl_logic_vector(31 downto 0);
        inclock         : in     vl_logic;
        wren            : in     vl_logic;
        q               : out    vl_logic_vector(31 downto 0)
    );
end RAM;
